// Code your testbench here
// or browse Examples
`include "top.sv"


